module orion_mem_ports
(
);

endmodule
