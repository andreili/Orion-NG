module orion
(
);

endmodule
