module orion_port_decoder
(
);

endmodule
